magic
tech sky130A
magscale 1 2
timestamp 1624412828
<< obsli1 >>
rect 1104 1785 184000 184977
<< obsm1 >>
rect 198 1640 184906 185008
<< metal2 >>
rect 754 186472 810 187272
rect 2318 186472 2374 187272
rect 3974 186472 4030 187272
rect 5538 186472 5594 187272
rect 7194 186472 7250 187272
rect 8850 186472 8906 187272
rect 10414 186472 10470 187272
rect 12070 186472 12126 187272
rect 13726 186472 13782 187272
rect 15290 186472 15346 187272
rect 16946 186472 17002 187272
rect 18602 186472 18658 187272
rect 20166 186472 20222 187272
rect 21822 186472 21878 187272
rect 23478 186472 23534 187272
rect 25042 186472 25098 187272
rect 26698 186472 26754 187272
rect 28354 186472 28410 187272
rect 29918 186472 29974 187272
rect 31574 186472 31630 187272
rect 33138 186472 33194 187272
rect 34794 186472 34850 187272
rect 36450 186472 36506 187272
rect 38014 186472 38070 187272
rect 39670 186472 39726 187272
rect 41326 186472 41382 187272
rect 42890 186472 42946 187272
rect 44546 186472 44602 187272
rect 46202 186472 46258 187272
rect 47766 186472 47822 187272
rect 49422 186472 49478 187272
rect 51078 186472 51134 187272
rect 52642 186472 52698 187272
rect 54298 186472 54354 187272
rect 55954 186472 56010 187272
rect 57518 186472 57574 187272
rect 59174 186472 59230 187272
rect 60830 186472 60886 187272
rect 62394 186472 62450 187272
rect 64050 186472 64106 187272
rect 65614 186472 65670 187272
rect 67270 186472 67326 187272
rect 68926 186472 68982 187272
rect 70490 186472 70546 187272
rect 72146 186472 72202 187272
rect 73802 186472 73858 187272
rect 75366 186472 75422 187272
rect 77022 186472 77078 187272
rect 78678 186472 78734 187272
rect 80242 186472 80298 187272
rect 81898 186472 81954 187272
rect 83554 186472 83610 187272
rect 85118 186472 85174 187272
rect 86774 186472 86830 187272
rect 88430 186472 88486 187272
rect 89994 186472 90050 187272
rect 91650 186472 91706 187272
rect 93306 186472 93362 187272
rect 94870 186472 94926 187272
rect 96526 186472 96582 187272
rect 98090 186472 98146 187272
rect 99746 186472 99802 187272
rect 101402 186472 101458 187272
rect 102966 186472 103022 187272
rect 104622 186472 104678 187272
rect 106278 186472 106334 187272
rect 107842 186472 107898 187272
rect 109498 186472 109554 187272
rect 111154 186472 111210 187272
rect 112718 186472 112774 187272
rect 114374 186472 114430 187272
rect 116030 186472 116086 187272
rect 117594 186472 117650 187272
rect 119250 186472 119306 187272
rect 120906 186472 120962 187272
rect 122470 186472 122526 187272
rect 124126 186472 124182 187272
rect 125690 186472 125746 187272
rect 127346 186472 127402 187272
rect 129002 186472 129058 187272
rect 130566 186472 130622 187272
rect 132222 186472 132278 187272
rect 133878 186472 133934 187272
rect 135442 186472 135498 187272
rect 137098 186472 137154 187272
rect 138754 186472 138810 187272
rect 140318 186472 140374 187272
rect 141974 186472 142030 187272
rect 143630 186472 143686 187272
rect 145194 186472 145250 187272
rect 146850 186472 146906 187272
rect 148506 186472 148562 187272
rect 150070 186472 150126 187272
rect 151726 186472 151782 187272
rect 153382 186472 153438 187272
rect 154946 186472 155002 187272
rect 156602 186472 156658 187272
rect 158166 186472 158222 187272
rect 159822 186472 159878 187272
rect 161478 186472 161534 187272
rect 163042 186472 163098 187272
rect 164698 186472 164754 187272
rect 166354 186472 166410 187272
rect 167918 186472 167974 187272
rect 169574 186472 169630 187272
rect 171230 186472 171286 187272
rect 172794 186472 172850 187272
rect 174450 186472 174506 187272
rect 176106 186472 176162 187272
rect 177670 186472 177726 187272
rect 179326 186472 179382 187272
rect 180982 186472 181038 187272
rect 182546 186472 182602 187272
rect 184202 186472 184258 187272
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88706 0 88762 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100482 0 100538 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131394 0 131450 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132866 0 132922 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152462 0 152518 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161110 0 161166 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163778 0 163834 800
rect 164146 0 164202 800
rect 164514 0 164570 800
rect 164882 0 164938 800
rect 165250 0 165306 800
rect 165618 0 165674 800
rect 166078 0 166134 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168286 0 168342 800
rect 168654 0 168710 800
rect 169022 0 169078 800
rect 169390 0 169446 800
rect 169758 0 169814 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176566 0 176622 800
rect 176934 0 176990 800
rect 177302 0 177358 800
rect 177762 0 177818 800
rect 178130 0 178186 800
rect 178498 0 178554 800
rect 178866 0 178922 800
rect 179234 0 179290 800
rect 179602 0 179658 800
rect 179970 0 180026 800
rect 180338 0 180394 800
rect 180706 0 180762 800
rect 181074 0 181130 800
rect 181534 0 181590 800
rect 181902 0 181958 800
rect 182270 0 182326 800
rect 182638 0 182694 800
rect 183006 0 183062 800
rect 183374 0 183430 800
rect 183742 0 183798 800
rect 184110 0 184166 800
rect 184478 0 184534 800
rect 184846 0 184902 800
<< obsm2 >>
rect 204 186416 698 186472
rect 866 186416 2262 186472
rect 2430 186416 3918 186472
rect 4086 186416 5482 186472
rect 5650 186416 7138 186472
rect 7306 186416 8794 186472
rect 8962 186416 10358 186472
rect 10526 186416 12014 186472
rect 12182 186416 13670 186472
rect 13838 186416 15234 186472
rect 15402 186416 16890 186472
rect 17058 186416 18546 186472
rect 18714 186416 20110 186472
rect 20278 186416 21766 186472
rect 21934 186416 23422 186472
rect 23590 186416 24986 186472
rect 25154 186416 26642 186472
rect 26810 186416 28298 186472
rect 28466 186416 29862 186472
rect 30030 186416 31518 186472
rect 31686 186416 33082 186472
rect 33250 186416 34738 186472
rect 34906 186416 36394 186472
rect 36562 186416 37958 186472
rect 38126 186416 39614 186472
rect 39782 186416 41270 186472
rect 41438 186416 42834 186472
rect 43002 186416 44490 186472
rect 44658 186416 46146 186472
rect 46314 186416 47710 186472
rect 47878 186416 49366 186472
rect 49534 186416 51022 186472
rect 51190 186416 52586 186472
rect 52754 186416 54242 186472
rect 54410 186416 55898 186472
rect 56066 186416 57462 186472
rect 57630 186416 59118 186472
rect 59286 186416 60774 186472
rect 60942 186416 62338 186472
rect 62506 186416 63994 186472
rect 64162 186416 65558 186472
rect 65726 186416 67214 186472
rect 67382 186416 68870 186472
rect 69038 186416 70434 186472
rect 70602 186416 72090 186472
rect 72258 186416 73746 186472
rect 73914 186416 75310 186472
rect 75478 186416 76966 186472
rect 77134 186416 78622 186472
rect 78790 186416 80186 186472
rect 80354 186416 81842 186472
rect 82010 186416 83498 186472
rect 83666 186416 85062 186472
rect 85230 186416 86718 186472
rect 86886 186416 88374 186472
rect 88542 186416 89938 186472
rect 90106 186416 91594 186472
rect 91762 186416 93250 186472
rect 93418 186416 94814 186472
rect 94982 186416 96470 186472
rect 96638 186416 98034 186472
rect 98202 186416 99690 186472
rect 99858 186416 101346 186472
rect 101514 186416 102910 186472
rect 103078 186416 104566 186472
rect 104734 186416 106222 186472
rect 106390 186416 107786 186472
rect 107954 186416 109442 186472
rect 109610 186416 111098 186472
rect 111266 186416 112662 186472
rect 112830 186416 114318 186472
rect 114486 186416 115974 186472
rect 116142 186416 117538 186472
rect 117706 186416 119194 186472
rect 119362 186416 120850 186472
rect 121018 186416 122414 186472
rect 122582 186416 124070 186472
rect 124238 186416 125634 186472
rect 125802 186416 127290 186472
rect 127458 186416 128946 186472
rect 129114 186416 130510 186472
rect 130678 186416 132166 186472
rect 132334 186416 133822 186472
rect 133990 186416 135386 186472
rect 135554 186416 137042 186472
rect 137210 186416 138698 186472
rect 138866 186416 140262 186472
rect 140430 186416 141918 186472
rect 142086 186416 143574 186472
rect 143742 186416 145138 186472
rect 145306 186416 146794 186472
rect 146962 186416 148450 186472
rect 148618 186416 150014 186472
rect 150182 186416 151670 186472
rect 151838 186416 153326 186472
rect 153494 186416 154890 186472
rect 155058 186416 156546 186472
rect 156714 186416 158110 186472
rect 158278 186416 159766 186472
rect 159934 186416 161422 186472
rect 161590 186416 162986 186472
rect 163154 186416 164642 186472
rect 164810 186416 166298 186472
rect 166466 186416 167862 186472
rect 168030 186416 169518 186472
rect 169686 186416 171174 186472
rect 171342 186416 172738 186472
rect 172906 186416 174394 186472
rect 174562 186416 176050 186472
rect 176218 186416 177614 186472
rect 177782 186416 179270 186472
rect 179438 186416 180926 186472
rect 181094 186416 182490 186472
rect 182658 186416 184146 186472
rect 184314 186416 184900 186472
rect 204 856 184900 186416
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1250 856
rect 1418 800 1618 856
rect 1786 800 1986 856
rect 2154 800 2354 856
rect 2522 800 2722 856
rect 2890 800 3090 856
rect 3258 800 3458 856
rect 3626 800 3826 856
rect 3994 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6862 856
rect 7030 800 7230 856
rect 7398 800 7598 856
rect 7766 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8794 856
rect 8962 800 9162 856
rect 9330 800 9530 856
rect 9698 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10634 856
rect 10802 800 11002 856
rect 11170 800 11370 856
rect 11538 800 11830 856
rect 11998 800 12198 856
rect 12366 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13302 856
rect 13470 800 13670 856
rect 13838 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15602 856
rect 15770 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16706 856
rect 16874 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17810 856
rect 17978 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19742 856
rect 19910 800 20110 856
rect 20278 800 20478 856
rect 20646 800 20846 856
rect 21014 800 21214 856
rect 21382 800 21582 856
rect 21750 800 21950 856
rect 22118 800 22318 856
rect 22486 800 22686 856
rect 22854 800 23054 856
rect 23222 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 26090 856
rect 26258 800 26458 856
rect 26626 800 26826 856
rect 26994 800 27286 856
rect 27454 800 27654 856
rect 27822 800 28022 856
rect 28190 800 28390 856
rect 28558 800 28758 856
rect 28926 800 29126 856
rect 29294 800 29494 856
rect 29662 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30598 856
rect 30766 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33634 856
rect 33802 800 34002 856
rect 34170 800 34370 856
rect 34538 800 34738 856
rect 34906 800 35198 856
rect 35366 800 35566 856
rect 35734 800 35934 856
rect 36102 800 36302 856
rect 36470 800 36670 856
rect 36838 800 37038 856
rect 37206 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38970 856
rect 39138 800 39338 856
rect 39506 800 39706 856
rect 39874 800 40074 856
rect 40242 800 40442 856
rect 40610 800 40810 856
rect 40978 800 41178 856
rect 41346 800 41546 856
rect 41714 800 41914 856
rect 42082 800 42282 856
rect 42450 800 42742 856
rect 42910 800 43110 856
rect 43278 800 43478 856
rect 43646 800 43846 856
rect 44014 800 44214 856
rect 44382 800 44582 856
rect 44750 800 44950 856
rect 45118 800 45318 856
rect 45486 800 45686 856
rect 45854 800 46054 856
rect 46222 800 46514 856
rect 46682 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47618 856
rect 47786 800 47986 856
rect 48154 800 48354 856
rect 48522 800 48722 856
rect 48890 800 49090 856
rect 49258 800 49458 856
rect 49626 800 49826 856
rect 49994 800 50286 856
rect 50454 800 50654 856
rect 50822 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51758 856
rect 51926 800 52126 856
rect 52294 800 52494 856
rect 52662 800 52862 856
rect 53030 800 53230 856
rect 53398 800 53598 856
rect 53766 800 53966 856
rect 54134 800 54426 856
rect 54594 800 54794 856
rect 54962 800 55162 856
rect 55330 800 55530 856
rect 55698 800 55898 856
rect 56066 800 56266 856
rect 56434 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57738 856
rect 57906 800 58198 856
rect 58366 800 58566 856
rect 58734 800 58934 856
rect 59102 800 59302 856
rect 59470 800 59670 856
rect 59838 800 60038 856
rect 60206 800 60406 856
rect 60574 800 60774 856
rect 60942 800 61142 856
rect 61310 800 61510 856
rect 61678 800 61970 856
rect 62138 800 62338 856
rect 62506 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63810 856
rect 63978 800 64178 856
rect 64346 800 64546 856
rect 64714 800 64914 856
rect 65082 800 65282 856
rect 65450 800 65742 856
rect 65910 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66846 856
rect 67014 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68318 856
rect 68486 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69422 856
rect 69590 800 69882 856
rect 70050 800 70250 856
rect 70418 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71354 856
rect 71522 800 71722 856
rect 71890 800 72090 856
rect 72258 800 72458 856
rect 72626 800 72826 856
rect 72994 800 73194 856
rect 73362 800 73654 856
rect 73822 800 74022 856
rect 74190 800 74390 856
rect 74558 800 74758 856
rect 74926 800 75126 856
rect 75294 800 75494 856
rect 75662 800 75862 856
rect 76030 800 76230 856
rect 76398 800 76598 856
rect 76766 800 76966 856
rect 77134 800 77426 856
rect 77594 800 77794 856
rect 77962 800 78162 856
rect 78330 800 78530 856
rect 78698 800 78898 856
rect 79066 800 79266 856
rect 79434 800 79634 856
rect 79802 800 80002 856
rect 80170 800 80370 856
rect 80538 800 80738 856
rect 80906 800 81198 856
rect 81366 800 81566 856
rect 81734 800 81934 856
rect 82102 800 82302 856
rect 82470 800 82670 856
rect 82838 800 83038 856
rect 83206 800 83406 856
rect 83574 800 83774 856
rect 83942 800 84142 856
rect 84310 800 84510 856
rect 84678 800 84878 856
rect 85046 800 85338 856
rect 85506 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88282 856
rect 88450 800 88650 856
rect 88818 800 89110 856
rect 89278 800 89478 856
rect 89646 800 89846 856
rect 90014 800 90214 856
rect 90382 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91686 856
rect 91854 800 92054 856
rect 92222 800 92422 856
rect 92590 800 92882 856
rect 93050 800 93250 856
rect 93418 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96194 856
rect 96362 800 96654 856
rect 96822 800 97022 856
rect 97190 800 97390 856
rect 97558 800 97758 856
rect 97926 800 98126 856
rect 98294 800 98494 856
rect 98662 800 98862 856
rect 99030 800 99230 856
rect 99398 800 99598 856
rect 99766 800 99966 856
rect 100134 800 100426 856
rect 100594 800 100794 856
rect 100962 800 101162 856
rect 101330 800 101530 856
rect 101698 800 101898 856
rect 102066 800 102266 856
rect 102434 800 102634 856
rect 102802 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104566 856
rect 104734 800 104934 856
rect 105102 800 105302 856
rect 105470 800 105670 856
rect 105838 800 106038 856
rect 106206 800 106406 856
rect 106574 800 106774 856
rect 106942 800 107142 856
rect 107310 800 107510 856
rect 107678 800 107878 856
rect 108046 800 108338 856
rect 108506 800 108706 856
rect 108874 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110546 856
rect 110714 800 110914 856
rect 111082 800 111282 856
rect 111450 800 111650 856
rect 111818 800 112110 856
rect 112278 800 112478 856
rect 112646 800 112846 856
rect 113014 800 113214 856
rect 113382 800 113582 856
rect 113750 800 113950 856
rect 114118 800 114318 856
rect 114486 800 114686 856
rect 114854 800 115054 856
rect 115222 800 115422 856
rect 115590 800 115882 856
rect 116050 800 116250 856
rect 116418 800 116618 856
rect 116786 800 116986 856
rect 117154 800 117354 856
rect 117522 800 117722 856
rect 117890 800 118090 856
rect 118258 800 118458 856
rect 118626 800 118826 856
rect 118994 800 119194 856
rect 119362 800 119562 856
rect 119730 800 120022 856
rect 120190 800 120390 856
rect 120558 800 120758 856
rect 120926 800 121126 856
rect 121294 800 121494 856
rect 121662 800 121862 856
rect 122030 800 122230 856
rect 122398 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123794 856
rect 123962 800 124162 856
rect 124330 800 124530 856
rect 124698 800 124898 856
rect 125066 800 125266 856
rect 125434 800 125634 856
rect 125802 800 126002 856
rect 126170 800 126370 856
rect 126538 800 126738 856
rect 126906 800 127106 856
rect 127274 800 127566 856
rect 127734 800 127934 856
rect 128102 800 128302 856
rect 128470 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130510 856
rect 130678 800 130878 856
rect 131046 800 131338 856
rect 131506 800 131706 856
rect 131874 800 132074 856
rect 132242 800 132442 856
rect 132610 800 132810 856
rect 132978 800 133178 856
rect 133346 800 133546 856
rect 133714 800 133914 856
rect 134082 800 134282 856
rect 134450 800 134650 856
rect 134818 800 135018 856
rect 135186 800 135478 856
rect 135646 800 135846 856
rect 136014 800 136214 856
rect 136382 800 136582 856
rect 136750 800 136950 856
rect 137118 800 137318 856
rect 137486 800 137686 856
rect 137854 800 138054 856
rect 138222 800 138422 856
rect 138590 800 138790 856
rect 138958 800 139250 856
rect 139418 800 139618 856
rect 139786 800 139986 856
rect 140154 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141090 856
rect 141258 800 141458 856
rect 141626 800 141826 856
rect 141994 800 142194 856
rect 142362 800 142562 856
rect 142730 800 143022 856
rect 143190 800 143390 856
rect 143558 800 143758 856
rect 143926 800 144126 856
rect 144294 800 144494 856
rect 144662 800 144862 856
rect 145030 800 145230 856
rect 145398 800 145598 856
rect 145766 800 145966 856
rect 146134 800 146334 856
rect 146502 800 146794 856
rect 146962 800 147162 856
rect 147330 800 147530 856
rect 147698 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 149002 856
rect 149170 800 149370 856
rect 149538 800 149738 856
rect 149906 800 150106 856
rect 150274 800 150566 856
rect 150734 800 150934 856
rect 151102 800 151302 856
rect 151470 800 151670 856
rect 151838 800 152038 856
rect 152206 800 152406 856
rect 152574 800 152774 856
rect 152942 800 153142 856
rect 153310 800 153510 856
rect 153678 800 153878 856
rect 154046 800 154246 856
rect 154414 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158478 856
rect 158646 800 158846 856
rect 159014 800 159214 856
rect 159382 800 159582 856
rect 159750 800 159950 856
rect 160118 800 160318 856
rect 160486 800 160686 856
rect 160854 800 161054 856
rect 161222 800 161422 856
rect 161590 800 161790 856
rect 161958 800 162250 856
rect 162418 800 162618 856
rect 162786 800 162986 856
rect 163154 800 163354 856
rect 163522 800 163722 856
rect 163890 800 164090 856
rect 164258 800 164458 856
rect 164626 800 164826 856
rect 164994 800 165194 856
rect 165362 800 165562 856
rect 165730 800 166022 856
rect 166190 800 166390 856
rect 166558 800 166758 856
rect 166926 800 167126 856
rect 167294 800 167494 856
rect 167662 800 167862 856
rect 168030 800 168230 856
rect 168398 800 168598 856
rect 168766 800 168966 856
rect 169134 800 169334 856
rect 169502 800 169702 856
rect 169870 800 170162 856
rect 170330 800 170530 856
rect 170698 800 170898 856
rect 171066 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173106 856
rect 173274 800 173474 856
rect 173642 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
rect 175574 800 175774 856
rect 175942 800 176142 856
rect 176310 800 176510 856
rect 176678 800 176878 856
rect 177046 800 177246 856
rect 177414 800 177706 856
rect 177874 800 178074 856
rect 178242 800 178442 856
rect 178610 800 178810 856
rect 178978 800 179178 856
rect 179346 800 179546 856
rect 179714 800 179914 856
rect 180082 800 180282 856
rect 180450 800 180650 856
rect 180818 800 181018 856
rect 181186 800 181478 856
rect 181646 800 181846 856
rect 182014 800 182214 856
rect 182382 800 182582 856
rect 182750 800 182950 856
rect 183118 800 183318 856
rect 183486 800 183686 856
rect 183854 800 184054 856
rect 184222 800 184422 856
rect 184590 800 184790 856
<< metal3 >>
rect 0 93576 800 93696
rect 184328 93576 185128 93696
<< obsm3 >>
rect 800 93776 184328 184993
rect 880 93496 184248 93776
rect 800 2143 184328 93496
<< metal4 >>
rect 4208 2128 4528 185008
rect 4868 2176 5188 184960
rect 5528 2176 5848 184960
rect 6188 2176 6508 184960
rect 19568 2128 19888 185008
rect 20228 2176 20548 184960
rect 20888 2176 21208 184960
rect 21548 2176 21868 184960
rect 34928 2128 35248 185008
rect 35588 2176 35908 184960
rect 36248 2176 36568 184960
rect 36908 2176 37228 184960
rect 50288 2128 50608 185008
rect 50948 2176 51268 184960
rect 51608 2176 51928 184960
rect 52268 2176 52588 184960
rect 65648 2128 65968 185008
rect 66308 2176 66628 184960
rect 66968 2176 67288 184960
rect 67628 2176 67948 184960
rect 81008 2128 81328 185008
rect 81668 2176 81988 184960
rect 82328 2176 82648 184960
rect 82988 2176 83308 184960
rect 96368 2128 96688 185008
rect 97028 2176 97348 184960
rect 97688 2176 98008 184960
rect 98348 2176 98668 184960
rect 111728 2128 112048 185008
rect 112388 2176 112708 184960
rect 113048 2176 113368 184960
rect 113708 2176 114028 184960
rect 127088 2128 127408 185008
rect 127748 2176 128068 184960
rect 128408 2176 128728 184960
rect 129068 2176 129388 184960
rect 142448 2128 142768 185008
rect 143108 2176 143428 184960
rect 143768 2176 144088 184960
rect 144428 2176 144748 184960
rect 157808 2128 158128 185008
rect 158468 2176 158788 184960
rect 159128 2176 159448 184960
rect 159788 2176 160108 184960
rect 173168 2128 173488 185008
rect 173828 2176 174148 184960
rect 174488 2176 174808 184960
rect 175148 2176 175468 184960
<< obsm4 >>
rect 15331 2483 19488 84693
rect 19968 2483 20148 84693
rect 20628 2483 20808 84693
rect 21288 2483 21468 84693
rect 21948 2483 34848 84693
rect 35328 2483 35508 84693
rect 35988 2483 36168 84693
rect 36648 2483 36828 84693
rect 37308 2483 50173 84693
<< labels >>
rlabel metal2 s 754 186472 810 187272 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 49422 186472 49478 187272 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 54298 186472 54354 187272 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 59174 186472 59230 187272 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 64050 186472 64106 187272 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 68926 186472 68982 187272 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 73802 186472 73858 187272 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 78678 186472 78734 187272 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 83554 186472 83610 187272 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 88430 186472 88486 187272 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 93306 186472 93362 187272 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5538 186472 5594 187272 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 98090 186472 98146 187272 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 102966 186472 103022 187272 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 107842 186472 107898 187272 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 112718 186472 112774 187272 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 117594 186472 117650 187272 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 122470 186472 122526 187272 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 127346 186472 127402 187272 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 132222 186472 132278 187272 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 137098 186472 137154 187272 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 141974 186472 142030 187272 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10414 186472 10470 187272 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 146850 186472 146906 187272 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 151726 186472 151782 187272 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 156602 186472 156658 187272 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 161478 186472 161534 187272 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 166354 186472 166410 187272 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 171230 186472 171286 187272 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 176106 186472 176162 187272 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 180982 186472 181038 187272 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15290 186472 15346 187272 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 20166 186472 20222 187272 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 25042 186472 25098 187272 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29918 186472 29974 187272 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 34794 186472 34850 187272 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 39670 186472 39726 187272 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 44546 186472 44602 187272 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 186472 2374 187272 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 51078 186472 51134 187272 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 55954 186472 56010 187272 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 60830 186472 60886 187272 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 65614 186472 65670 187272 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 70490 186472 70546 187272 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 75366 186472 75422 187272 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 80242 186472 80298 187272 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 85118 186472 85174 187272 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 89994 186472 90050 187272 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 94870 186472 94926 187272 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7194 186472 7250 187272 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 99746 186472 99802 187272 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 104622 186472 104678 187272 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 109498 186472 109554 187272 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 114374 186472 114430 187272 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 119250 186472 119306 187272 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 124126 186472 124182 187272 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 129002 186472 129058 187272 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 133878 186472 133934 187272 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 138754 186472 138810 187272 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 143630 186472 143686 187272 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12070 186472 12126 187272 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 148506 186472 148562 187272 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 153382 186472 153438 187272 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 158166 186472 158222 187272 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 163042 186472 163098 187272 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 167918 186472 167974 187272 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 172794 186472 172850 187272 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 177670 186472 177726 187272 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 182546 186472 182602 187272 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16946 186472 17002 187272 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21822 186472 21878 187272 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26698 186472 26754 187272 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 31574 186472 31630 187272 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 36450 186472 36506 187272 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 41326 186472 41382 187272 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 46202 186472 46258 187272 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3974 186472 4030 187272 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 52642 186472 52698 187272 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 57518 186472 57574 187272 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 62394 186472 62450 187272 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 67270 186472 67326 187272 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 72146 186472 72202 187272 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 77022 186472 77078 187272 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 81898 186472 81954 187272 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 86774 186472 86830 187272 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 91650 186472 91706 187272 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 96526 186472 96582 187272 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8850 186472 8906 187272 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 101402 186472 101458 187272 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 106278 186472 106334 187272 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 111154 186472 111210 187272 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 116030 186472 116086 187272 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 120906 186472 120962 187272 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 125690 186472 125746 187272 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 130566 186472 130622 187272 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 135442 186472 135498 187272 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 140318 186472 140374 187272 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 145194 186472 145250 187272 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13726 186472 13782 187272 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 150070 186472 150126 187272 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 154946 186472 155002 187272 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 159822 186472 159878 187272 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 164698 186472 164754 187272 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 169574 186472 169630 187272 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 174450 186472 174506 187272 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 179326 186472 179382 187272 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 184202 186472 184258 187272 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18602 186472 18658 187272 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 23478 186472 23534 187272 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 28354 186472 28410 187272 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 33138 186472 33194 187272 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 38014 186472 38070 187272 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42890 186472 42946 187272 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 47766 186472 47822 187272 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 184328 93576 185128 93696 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 168286 0 168342 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 183006 0 183062 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 185008 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 185008 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 185008 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 185008 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 185008 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 185008 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 185008 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 185008 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 185008 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 185008 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 185008 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 185008 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 184960 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 184960 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 184960 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 184960 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 184960 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 184960 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 184960 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 184960 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 184960 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 184960 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 184960 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 184960 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 184960 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 184960 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 184960 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 184960 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 184960 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 184960 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 184960 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 184960 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 184960 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 184960 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 184960 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 184960 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 184960 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 184960 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 184960 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 184960 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 184960 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 184960 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 184960 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 184960 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 184960 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 184960 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 184960 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 184960 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 185128 187272
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 52614182
string GDS_START 1407294
<< end >>

